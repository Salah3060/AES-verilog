

module invShiftRow_tb() ;

reg [0:127] data ;
wire[0:127] out;

invShiftRow INV(data , out);

initial
 begin
    data = 128'h_00_00_00; #100;
    data = 128'h6353e08c0960e104cd70b751bacad0e7; 
    $monitor("--> out %h" , out);  

end 





endmodule